localparam[15:0] DATAI_REG_ADDR = 16'h0000;
localparam[15:0] DATAO_REG_ADDR = 16'h0004;
localparam[15:0] DIR_REG_ADDR = 16'h0008;
localparam[15:0] ICR_REG_ADDR = 16'h0f00;
localparam[15:0] RIS_REG_ADDR = 16'h0f04;
localparam[15:0] IM_REG_ADDR = 16'h0f08;
localparam[15:0] MIS_REG_ADDR = 16'h0f0c;

localparam  GPIO8_DATAI_REG_DATAI = 0,
            GPIO8_DATAI_REG_DATAI_LEN = 8,
            GPIO8_DATAO_REG_DATAO = 0,
            GPIO8_DATAO_REG_DATAO_LEN = 8,
            GPIO8_DIR_REG_DIR = 0,
            GPIO8_DIR_REG_DIR_LEN = 8,
            GPIO8_PIN0_HI_FLAG = 32'h1,
            GPIO8_PIN1_HI_FLAG = 32'h2,
            GPIO8_PIN2_HI_FLAG = 32'h4,
            GPIO8_PIN3_HI_FLAG = 32'h8,
            GPIO8_PIN4_HI_FLAG = 32'h10,
            GPIO8_PIN5_HI_FLAG = 32'h20,
            GPIO8_PIN6_HI_FLAG = 32'h40,
            GPIO8_PIN7_HI_FLAG = 32'h80,
            GPIO8_PIN0_LO_FLAG = 32'h100,
            GPIO8_PIN1_LO_FLAG = 32'h200,
            GPIO8_PIN2_LO_FLAG = 32'h400,
            GPIO8_PIN3_LO_FLAG = 32'h800,
            GPIO8_PIN4_LO_FLAG = 32'h1000,
            GPIO8_PIN5_LO_FLAG = 32'h2000,
            GPIO8_PIN6_LO_FLAG = 32'h4000,
            GPIO8_PIN7_LO_FLAG = 32'h8000,
            GPIO8_PIN0_PE_FLAG = 32'h10000,
            GPIO8_PIN1_PE_FLAG = 32'h20000,
            GPIO8_PIN2_PE_FLAG = 32'h40000,
            GPIO8_PIN3_PE_FLAG = 32'h80000,
            GPIO8_PIN4_PE_FLAG = 32'h100000,
            GPIO8_PIN5_PE_FLAG = 32'h200000,
            GPIO8_PIN6_PE_FLAG = 32'h400000,
            GPIO8_PIN7_PE_FLAG = 32'h800000,
            GPIO8_PIN0_NE_FLAG = 32'h1000000,
            GPIO8_PIN1_NE_FLAG = 32'h2000000,
            GPIO8_PIN2_NE_FLAG = 32'h4000000,
            GPIO8_PIN3_NE_FLAG = 32'h8000000,
            GPIO8_PIN4_NE_FLAG = 32'h10000000,
            GPIO8_PIN5_NE_FLAG = 32'h20000000,
            GPIO8_PIN6_NE_FLAG = 32'h40000000,
            GPIO8_PIN7_NE_FLAG = 32'h80000000;
